interface intf();
  logic[7:0] A,B;
  logic[3:0] ALU_Sel;
  logic [7:0] ALU_Out;
  logic CarryOut;
endinterface